`define ADPLL_ADDR_W 5

`define ALPHA_L (`ADPLL_ADDR_W'd0)
`define ALPHA_M (`ADPLL_ADDR_W'd1)
`define ALPHA_S_RX (`ADPLL_ADDR_W'd2)
`define ALPHA_S_TX (`ADPLL_ADDR_W'd3)
`define BETA (`ADPLL_ADDR_W'd4)
`define LAMBDA_RX (`ADPLL_ADDR_W'd5)
`define LAMBDA_TX (`ADPLL_ADDR_W'd6)
`define IIR_N_RX (`ADPLL_ADDR_W'd7)
`define IIR_N_TX (`ADPLL_ADDR_W'd8)
`define FCW_MOD (`ADPLL_ADDR_W'd9)
`define DCO_C_L_WORD_TEST (`ADPLL_ADDR_W'd10)
`define DCO_C_M_WORD_TEST (`ADPLL_ADDR_W'd11)
`define DCO_C_S_WORD_TEST (`ADPLL_ADDR_W'd12)
`define DCO_PD_TEST (`ADPLL_ADDR_W'd13)
`define TDC_PD_TEST (`ADPLL_ADDR_W'd14)
`define TDC_PD_INJ_TEST (`ADPLL_ADDR_W'd15)
`define TDC_CTR_FREQ (`ADPLL_ADDR_W'd16)
`define DCO_OSC_GAIN (`ADPLL_ADDR_W'd17)
`define ADPLL_SOFT_RST (`ADPLL_ADDR_W'd18)
