// Created by ihdl
`timescale 10ps/1ps

`celldefine

module XNR3EHD(O, I1, I2, I3);
   output O;
   input I1, I2, I3;

//Function Block
`protect
   xnor g1(O, I1, I2, I3);

//Specify Block
   specify

      //  Module Path Delay (state dependent)
      if (I1 == 0 && I2 == 1) (I3 *> O) = (6.00:6.00:6.00, 5.94:5.94:5.94);
      if (I1 == 1 && I2 == 1) (I3 *> O) = (7.42:7.42:7.42, 5.85:5.85:5.85);
      if (I1 == 0 && I2 == 0) (I3 *> O) = (7.34:7.34:7.34, 5.91:5.91:5.91);
      if (I1 == 1 && I2 == 0) (I3 *> O) = (6.05:6.05:6.05, 5.90:5.90:5.90);
      ifnone (I3 *> O) = (6.05:6.05:6.05, 5.90:5.90:5.90);
      if (I1 == 0 && I3 == 0) (I2 *> O) = (11.19:11.19:11.19, 9.35:9.35:9.35);
      if (I1 == 1 && I3 == 0) (I2 *> O) = (9.69:9.69:9.69, 9.82:9.82:9.82);
      if (I1 == 0 && I3 == 1) (I2 *> O) = (9.55:9.55:9.55, 10.19:10.19:10.19);
      if (I1 == 1 && I3 == 1) (I2 *> O) = (11.26:11.26:11.26, 9.05:9.05:9.05);
      ifnone (I2 *> O) = (11.26:11.26:11.26, 9.05:9.05:9.05);
      if (I2 == 0 && I3 == 0) (I1 *> O) = (17.15:17.15:17.15, 14.30:14.30:14.30);
      if (I2 == 1 && I3 == 0) (I1 *> O) = (12.16:12.16:12.16, 12.56:12.56:12.56);
      if (I2 == 0 && I3 == 1) (I1 *> O) = (12.12:12.12:12.12, 12.54:12.54:12.54);
      if (I2 == 1 && I3 == 1) (I1 *> O) = (17.04:17.04:17.04, 14.39:14.39:14.39);
      ifnone (I1 *> O) = (17.04:17.04:17.04, 14.39:14.39:14.39);

      //  Module Path Delay
   endspecify
`endprotect
endmodule

`endcelldefine
