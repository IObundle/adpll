// Created by ihdl
`timescale 10ps/1ps

`celldefine

module AO2222EHD(O, A1, A2, B1, B2, C1, C2, D1, D2);
   output O;
   input A1, A2, B1, B2, C1, C2, D1, D2;

//Function Block
`protect
   and g1(o1, B1, B2);
   and g3(o2, A1, A2);
   and g4(o3, C1, C2);
   and g5(o4, D1, D2);
   nor g2(o5, o1, o2, o3, o4);
   not g6(O,o5);

//Specify Block
   specify

      //  Module Path Delay (state dependent)
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 0 && C1 == 0 && C2 == 1) (D1 *> O) = (5.70:5.70:5.70, 6.63:6.63:6.63);
      if (A1 == 1 && A2 == 0 && B1 == 1 && B2 == 0 && C1 == 1 && C2 == 0) (D1 *> O) = (6.22:6.22:6.22, 8.01:8.01:8.01);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 1 && C1 == 0 && C2 == 0) (D1 *> O) = (5.69:5.69:5.69, 5.52:5.52:5.52);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 0 && C1 == 0 && C2 == 0) (D1 *> O) = (5.69:5.69:5.69, 5.52:5.52:5.52);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 1 && C1 == 0 && C2 == 1) (D1 *> O) = (5.70:5.70:5.70, 6.63:6.63:6.63);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 0 && C1 == 0 && C2 == 1) (D1 *> O) = (5.70:5.70:5.70, 6.63:6.63:6.63);
      if (A1 == 1 && A2 == 0 && B1 == 1 && B2 == 0 && C1 == 0 && C2 == 0) (D1 *> O) = (5.69:5.69:5.69, 5.52:5.52:5.52);
      if (A1 == 1 && A2 == 0 && B1 == 1 && B2 == 0 && C1 == 0 && C2 == 1) (D1 *> O) = (5.70:5.70:5.70, 6.63:6.63:6.63);
      if (A1 == 0 && A2 == 1 && B1 == 1 && B2 == 0 && C1 == 1 && C2 == 0) (D1 *> O) = (6.22:6.22:6.22, 8.01:8.01:8.01);
      if (A1 == 0 && A2 == 0 && B1 == 1 && B2 == 0 && C1 == 1 && C2 == 0) (D1 *> O) = (6.22:6.22:6.22, 8.01:8.01:8.01);
      if (A1 == 0 && A2 == 1 && B1 == 1 && B2 == 0 && C1 == 0 && C2 == 0) (D1 *> O) = (5.69:5.69:5.69, 5.52:5.52:5.52);
      if (A1 == 0 && A2 == 1 && B1 == 1 && B2 == 0 && C1 == 0 && C2 == 1) (D1 *> O) = (5.70:5.70:5.70, 6.63:6.63:6.63);
      if (A1 == 0 && A2 == 0 && B1 == 1 && B2 == 0 && C1 == 0 && C2 == 0) (D1 *> O) = (5.69:5.69:5.69, 5.52:5.52:5.52);
      if (A1 == 0 && A2 == 0 && B1 == 1 && B2 == 0 && C1 == 0 && C2 == 1) (D1 *> O) = (5.70:5.70:5.70, 6.63:6.63:6.63);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 1 && C1 == 1 && C2 == 0) (D1 *> O) = (6.22:6.22:6.22, 8.01:8.01:8.01);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 0 && C1 == 1 && C2 == 0) (D1 *> O) = (6.22:6.22:6.22, 8.01:8.01:8.01);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 1 && C1 == 0 && C2 == 0) (D1 *> O) = (5.69:5.69:5.69, 5.52:5.52:5.52);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 0 && C1 == 0 && C2 == 0) (D1 *> O) = (5.69:5.69:5.69, 5.52:5.52:5.52);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 1 && C1 == 0 && C2 == 1) (D1 *> O) = (5.70:5.70:5.70, 6.63:6.63:6.63);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 1 && C1 == 1 && C2 == 0) (D1 *> O) = (6.22:6.22:6.22, 8.01:8.01:8.01);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 0 && C1 == 0 && C2 == 1) (D1 *> O) = (5.70:5.70:5.70, 6.63:6.63:6.63);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 0 && C1 == 1 && C2 == 0) (D1 *> O) = (6.22:6.22:6.22, 8.01:8.01:8.01);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 1 && C1 == 1 && C2 == 0) (D1 *> O) = (6.22:6.22:6.22, 8.01:8.01:8.01);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 0 && C1 == 1 && C2 == 0) (D1 *> O) = (6.23:6.23:6.23, 8.01:8.01:8.01);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 1 && C1 == 0 && C2 == 0) (D1 *> O) = (5.69:5.69:5.69, 5.52:5.52:5.52);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 0 && C1 == 0 && C2 == 0) (D1 *> O) = (5.69:5.69:5.69, 5.52:5.52:5.52);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 1 && C1 == 0 && C2 == 1) (D1 *> O) = (5.70:5.70:5.70, 6.63:6.63:6.63);
      ifnone (D1 *> O) = (5.70:5.70:5.70, 6.63:6.63:6.63);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 1 && C1 == 1 && C2 == 0) (D2 *> O) = (6.29:6.29:6.29, 8.66:8.66:8.66);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 0 && C1 == 1 && C2 == 0) (D2 *> O) = (6.29:6.29:6.29, 8.66:8.66:8.66);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 1 && C1 == 0 && C2 == 0) (D2 *> O) = (5.77:5.77:5.77, 6.04:6.04:6.04);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 0 && C1 == 0 && C2 == 0) (D2 *> O) = (5.77:5.77:5.77, 6.04:6.04:6.04);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 1 && C1 == 1 && C2 == 0) (D2 *> O) = (6.29:6.29:6.29, 8.66:8.66:8.66);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 1 && C1 == 0 && C2 == 1) (D2 *> O) = (5.78:5.78:5.78, 7.31:7.31:7.31);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 0 && C1 == 0 && C2 == 1) (D2 *> O) = (5.78:5.78:5.78, 7.31:7.31:7.31);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 0 && C1 == 1 && C2 == 0) (D2 *> O) = (6.29:6.29:6.29, 8.66:8.66:8.66);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 1 && C1 == 1 && C2 == 0) (D2 *> O) = (6.29:6.29:6.29, 8.66:8.66:8.66);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 0 && C1 == 1 && C2 == 0) (D2 *> O) = (6.29:6.29:6.29, 8.66:8.66:8.66);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 1 && C1 == 0 && C2 == 0) (D2 *> O) = (5.77:5.77:5.77, 6.04:6.04:6.04);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 0 && C1 == 0 && C2 == 0) (D2 *> O) = (5.77:5.77:5.77, 6.04:6.04:6.04);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 1 && C1 == 0 && C2 == 1) (D2 *> O) = (5.78:5.78:5.78, 7.31:7.31:7.31);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 0 && C1 == 0 && C2 == 1) (D2 *> O) = (5.78:5.78:5.78, 7.31:7.31:7.31);
      if (A1 == 1 && A2 == 0 && B1 == 1 && B2 == 0 && C1 == 1 && C2 == 0) (D2 *> O) = (6.29:6.29:6.29, 8.66:8.66:8.66);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 1 && C1 == 0 && C2 == 0) (D2 *> O) = (5.77:5.77:5.77, 6.04:6.04:6.04);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 0 && C1 == 0 && C2 == 0) (D2 *> O) = (5.77:5.77:5.77, 6.04:6.04:6.04);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 1 && C1 == 0 && C2 == 1) (D2 *> O) = (5.78:5.78:5.78, 7.31:7.31:7.31);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 0 && C1 == 0 && C2 == 1) (D2 *> O) = (5.78:5.78:5.78, 7.31:7.31:7.31);
      if (A1 == 1 && A2 == 0 && B1 == 1 && B2 == 0 && C1 == 0 && C2 == 0) (D2 *> O) = (5.77:5.77:5.77, 6.04:6.04:6.04);
      if (A1 == 0 && A2 == 1 && B1 == 1 && B2 == 0 && C1 == 1 && C2 == 0) (D2 *> O) = (6.29:6.29:6.29, 8.66:8.66:8.66);
      if (A1 == 1 && A2 == 0 && B1 == 1 && B2 == 0 && C1 == 0 && C2 == 1) (D2 *> O) = (5.78:5.78:5.78, 7.31:7.31:7.31);
      if (A1 == 0 && A2 == 0 && B1 == 1 && B2 == 0 && C1 == 1 && C2 == 0) (D2 *> O) = (6.29:6.29:6.29, 8.66:8.66:8.66);
      if (A1 == 0 && A2 == 1 && B1 == 1 && B2 == 0 && C1 == 0 && C2 == 0) (D2 *> O) = (5.77:5.77:5.77, 6.04:6.04:6.04);
      if (A1 == 0 && A2 == 1 && B1 == 1 && B2 == 0 && C1 == 0 && C2 == 1) (D2 *> O) = (5.78:5.78:5.78, 7.31:7.31:7.31);
      if (A1 == 0 && A2 == 0 && B1 == 1 && B2 == 0 && C1 == 0 && C2 == 0) (D2 *> O) = (5.77:5.77:5.77, 6.04:6.04:6.04);
      if (A1 == 0 && A2 == 0 && B1 == 1 && B2 == 0 && C1 == 0 && C2 == 1) (D2 *> O) = (5.78:5.78:5.78, 7.31:7.31:7.31);
      ifnone (D2 *> O) = (5.78:5.78:5.78, 7.31:7.31:7.31);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 0 && D1 == 0 && D2 == 0) (C1 *> O) = (6.85:6.85:6.85, 7.10:7.10:7.10);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 1 && D1 == 0 && D2 == 1) (C1 *> O) = (6.52:6.52:6.52, 8.31:8.31:8.31);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 0 && D1 == 0 && D2 == 1) (C1 *> O) = (6.52:6.52:6.52, 8.31:8.31:8.31);
      if (A1 == 1 && A2 == 0 && B1 == 1 && B2 == 0 && D1 == 1 && D2 == 0) (C1 *> O) = (6.83:6.83:6.83, 9.13:9.13:9.13);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 1 && D1 == 0 && D2 == 0) (C1 *> O) = (6.85:6.85:6.85, 7.10:7.10:7.10);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 0 && D1 == 0 && D2 == 0) (C1 *> O) = (6.85:6.85:6.85, 7.10:7.10:7.10);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 1 && D1 == 0 && D2 == 1) (C1 *> O) = (6.52:6.52:6.52, 8.31:8.31:8.31);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 0 && D1 == 0 && D2 == 1) (C1 *> O) = (6.52:6.52:6.52, 8.31:8.31:8.31);
      if (A1 == 1 && A2 == 0 && B1 == 1 && B2 == 0 && D1 == 0 && D2 == 0) (C1 *> O) = (6.84:6.84:6.84, 7.10:7.10:7.10);
      if (A1 == 0 && A2 == 1 && B1 == 1 && B2 == 0 && D1 == 1 && D2 == 0) (C1 *> O) = (6.83:6.83:6.83, 9.13:9.13:9.13);
      if (A1 == 1 && A2 == 0 && B1 == 1 && B2 == 0 && D1 == 0 && D2 == 1) (C1 *> O) = (6.52:6.52:6.52, 8.31:8.31:8.31);
      if (A1 == 0 && A2 == 0 && B1 == 1 && B2 == 0 && D1 == 1 && D2 == 0) (C1 *> O) = (6.83:6.83:6.83, 9.13:9.13:9.13);
      if (A1 == 0 && A2 == 1 && B1 == 1 && B2 == 0 && D1 == 0 && D2 == 0) (C1 *> O) = (6.84:6.84:6.84, 7.10:7.10:7.10);
      if (A1 == 0 && A2 == 1 && B1 == 1 && B2 == 0 && D1 == 0 && D2 == 1) (C1 *> O) = (6.52:6.52:6.52, 8.31:8.31:8.31);
      if (A1 == 0 && A2 == 0 && B1 == 1 && B2 == 0 && D1 == 0 && D2 == 0) (C1 *> O) = (6.85:6.85:6.85, 7.10:7.10:7.10);
      if (A1 == 0 && A2 == 0 && B1 == 1 && B2 == 0 && D1 == 0 && D2 == 1) (C1 *> O) = (6.52:6.52:6.52, 8.31:8.31:8.31);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 1 && D1 == 1 && D2 == 0) (C1 *> O) = (6.83:6.83:6.83, 9.13:9.13:9.13);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 0 && D1 == 1 && D2 == 0) (C1 *> O) = (6.83:6.83:6.83, 9.13:9.13:9.13);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 1 && D1 == 0 && D2 == 0) (C1 *> O) = (6.84:6.84:6.84, 7.10:7.10:7.10);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 0 && D1 == 0 && D2 == 0) (C1 *> O) = (6.85:6.85:6.85, 7.10:7.10:7.10);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 1 && D1 == 1 && D2 == 0) (C1 *> O) = (6.83:6.83:6.83, 9.13:9.13:9.13);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 1 && D1 == 0 && D2 == 1) (C1 *> O) = (6.52:6.52:6.52, 8.31:8.31:8.31);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 0 && D1 == 1 && D2 == 0) (C1 *> O) = (6.83:6.83:6.83, 9.13:9.13:9.13);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 0 && D1 == 0 && D2 == 1) (C1 *> O) = (6.52:6.52:6.52, 8.31:8.31:8.31);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 1 && D1 == 1 && D2 == 0) (C1 *> O) = (6.83:6.83:6.83, 9.13:9.13:9.13);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 0 && D1 == 1 && D2 == 0) (C1 *> O) = (6.83:6.83:6.83, 9.13:9.13:9.13);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 1 && D1 == 0 && D2 == 0) (C1 *> O) = (6.84:6.84:6.84, 7.10:7.10:7.10);
      ifnone (C1 *> O) = (6.84:6.84:6.84, 7.10:7.10:7.10);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 1 && D1 == 1 && D2 == 0) (C2 *> O) = (7.15:7.15:7.15, 10.34:10.34:10.34);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 0 && D1 == 1 && D2 == 0) (C2 *> O) = (7.15:7.15:7.15, 10.34:10.34:10.34);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 1 && D1 == 0 && D2 == 0) (C2 *> O) = (7.17:7.17:7.17, 8.06:8.06:8.06);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 0 && D1 == 0 && D2 == 0) (C2 *> O) = (7.17:7.17:7.17, 8.06:8.06:8.06);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 1 && D1 == 1 && D2 == 0) (C2 *> O) = (7.15:7.15:7.15, 10.34:10.34:10.34);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 1 && D1 == 0 && D2 == 1) (C2 *> O) = (6.84:6.84:6.84, 9.55:9.55:9.55);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 0 && D1 == 1 && D2 == 0) (C2 *> O) = (7.15:7.15:7.15, 10.34:10.34:10.34);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 0 && D1 == 0 && D2 == 1) (C2 *> O) = (6.84:6.84:6.84, 9.55:9.55:9.55);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 1 && D1 == 1 && D2 == 0) (C2 *> O) = (7.15:7.15:7.15, 10.34:10.34:10.34);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 0 && D1 == 1 && D2 == 0) (C2 *> O) = (7.15:7.15:7.15, 10.34:10.34:10.34);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 1 && D1 == 0 && D2 == 0) (C2 *> O) = (7.17:7.17:7.17, 8.06:8.06:8.06);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 0 && D1 == 0 && D2 == 0) (C2 *> O) = (7.17:7.17:7.17, 8.06:8.06:8.06);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 1 && D1 == 0 && D2 == 1) (C2 *> O) = (6.84:6.84:6.84, 9.55:9.55:9.55);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 0 && D1 == 0 && D2 == 1) (C2 *> O) = (6.84:6.84:6.84, 9.55:9.55:9.55);
      if (A1 == 1 && A2 == 0 && B1 == 1 && B2 == 0 && D1 == 1 && D2 == 0) (C2 *> O) = (7.15:7.15:7.15, 10.34:10.34:10.34);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 1 && D1 == 0 && D2 == 0) (C2 *> O) = (7.17:7.17:7.17, 8.06:8.06:8.06);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 0 && D1 == 0 && D2 == 0) (C2 *> O) = (7.17:7.17:7.17, 8.06:8.06:8.06);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 1 && D1 == 0 && D2 == 1) (C2 *> O) = (6.84:6.84:6.84, 9.55:9.55:9.55);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 0 && D1 == 0 && D2 == 1) (C2 *> O) = (6.84:6.84:6.84, 9.55:9.55:9.55);
      if (A1 == 1 && A2 == 0 && B1 == 1 && B2 == 0 && D1 == 0 && D2 == 0) (C2 *> O) = (7.17:7.17:7.17, 8.06:8.06:8.06);
      if (A1 == 0 && A2 == 1 && B1 == 1 && B2 == 0 && D1 == 1 && D2 == 0) (C2 *> O) = (7.15:7.15:7.15, 10.34:10.34:10.34);
      if (A1 == 1 && A2 == 0 && B1 == 1 && B2 == 0 && D1 == 0 && D2 == 1) (C2 *> O) = (6.84:6.84:6.84, 9.55:9.55:9.55);
      if (A1 == 0 && A2 == 0 && B1 == 1 && B2 == 0 && D1 == 1 && D2 == 0) (C2 *> O) = (7.15:7.15:7.15, 10.34:10.34:10.34);
      if (A1 == 0 && A2 == 1 && B1 == 1 && B2 == 0 && D1 == 0 && D2 == 0) (C2 *> O) = (7.17:7.17:7.17, 8.06:8.06:8.06);
      if (A1 == 0 && A2 == 1 && B1 == 1 && B2 == 0 && D1 == 0 && D2 == 1) (C2 *> O) = (6.84:6.84:6.84, 9.55:9.55:9.55);
      if (A1 == 0 && A2 == 0 && B1 == 1 && B2 == 0 && D1 == 0 && D2 == 0) (C2 *> O) = (7.17:7.17:7.17, 8.06:8.06:8.06);
      if (A1 == 0 && A2 == 0 && B1 == 1 && B2 == 0 && D1 == 0 && D2 == 1) (C2 *> O) = (6.84:6.84:6.84, 9.55:9.55:9.55);
      ifnone (C2 *> O) = (6.84:6.84:6.84, 9.55:9.55:9.55);
      if (A1 == 1 && A2 == 0 && C1 == 0 && C2 == 1 && D1 == 1 && D2 == 0) (B1 *> O) = (7.22:7.22:7.22, 8.38:8.38:8.38);
      if (A1 == 1 && A2 == 0 && C1 == 0 && C2 == 0 && D1 == 1 && D2 == 0) (B1 *> O) = (7.23:7.23:7.23, 8.38:8.38:8.38);
      if (A1 == 1 && A2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 0) (B1 *> O) = (7.24:7.24:7.24, 8.37:8.37:8.37);
      if (A1 == 1 && A2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 0) (B1 *> O) = (7.25:7.25:7.25, 8.37:8.37:8.37);
      if (A1 == 0 && A2 == 1 && C1 == 0 && C2 == 1 && D1 == 1 && D2 == 0) (B1 *> O) = (6.67:6.67:6.67, 7.08:7.08:7.08);
      if (A1 == 1 && A2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 1) (B1 *> O) = (7.22:7.22:7.22, 8.38:8.38:8.38);
      if (A1 == 0 && A2 == 1 && C1 == 0 && C2 == 0 && D1 == 1 && D2 == 0) (B1 *> O) = (6.68:6.68:6.68, 7.08:7.08:7.08);
      if (A1 == 1 && A2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 1) (B1 *> O) = (7.23:7.23:7.23, 8.38:8.38:8.38);
      if (A1 == 0 && A2 == 0 && C1 == 0 && C2 == 1 && D1 == 1 && D2 == 0) (B1 *> O) = (6.66:6.66:6.66, 5.92:5.92:5.92);
      if (A1 == 0 && A2 == 0 && C1 == 0 && C2 == 0 && D1 == 1 && D2 == 0) (B1 *> O) = (6.67:6.67:6.67, 5.92:5.92:5.92);
      if (A1 == 0 && A2 == 1 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 0) (B1 *> O) = (6.69:6.69:6.69, 7.07:7.07:7.07);
      if (A1 == 0 && A2 == 1 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 0) (B1 *> O) = (6.71:6.71:6.71, 7.07:7.07:7.07);
      if (A1 == 0 && A2 == 1 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 1) (B1 *> O) = (6.67:6.67:6.67, 7.08:7.08:7.08);
      if (A1 == 0 && A2 == 1 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 1) (B1 *> O) = (6.68:6.68:6.68, 7.08:7.08:7.08);
      if (A1 == 1 && A2 == 0 && C1 == 1 && C2 == 0 && D1 == 1 && D2 == 0) (B1 *> O) = (7.22:7.22:7.22, 8.38:8.38:8.38);
      if (A1 == 0 && A2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 0) (B1 *> O) = (6.68:6.68:6.68, 5.91:5.91:5.91);
      if (A1 == 0 && A2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 0) (B1 *> O) = (6.70:6.70:6.70, 5.91:5.91:5.91);
      if (A1 == 0 && A2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 1) (B1 *> O) = (6.66:6.66:6.66, 5.92:5.92:5.92);
      if (A1 == 0 && A2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 1) (B1 *> O) = (6.67:6.67:6.67, 5.92:5.92:5.92);
      if (A1 == 1 && A2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 0) (B1 *> O) = (7.24:7.24:7.24, 8.37:8.37:8.37);
      if (A1 == 0 && A2 == 1 && C1 == 1 && C2 == 0 && D1 == 1 && D2 == 0) (B1 *> O) = (6.67:6.67:6.67, 7.08:7.08:7.08);
      if (A1 == 1 && A2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 1) (B1 *> O) = (7.22:7.22:7.22, 8.38:8.38:8.38);
      if (A1 == 0 && A2 == 0 && C1 == 1 && C2 == 0 && D1 == 1 && D2 == 0) (B1 *> O) = (6.66:6.66:6.66, 5.92:5.92:5.92);
      if (A1 == 0 && A2 == 1 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 0) (B1 *> O) = (6.69:6.69:6.69, 7.07:7.07:7.07);
      if (A1 == 0 && A2 == 1 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 1) (B1 *> O) = (6.67:6.67:6.67, 7.08:7.08:7.08);
      if (A1 == 0 && A2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 0) (B1 *> O) = (6.68:6.68:6.68, 5.91:5.91:5.91);
      if (A1 == 0 && A2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 1) (B1 *> O) = (6.66:6.66:6.66, 5.92:5.92:5.92);
      ifnone (B1 *> O) = (6.66:6.66:6.66, 5.92:5.92:5.92);
      if (A1 == 0 && A2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 1) (B2 *> O) = (6.74:6.74:6.74, 6.43:6.43:6.43);
      if (A1 == 1 && A2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 0) (B2 *> O) = (7.31:7.31:7.31, 9.02:9.02:9.02);
      if (A1 == 0 && A2 == 1 && C1 == 1 && C2 == 0 && D1 == 1 && D2 == 0) (B2 *> O) = (6.74:6.74:6.74, 7.75:7.75:7.75);
      if (A1 == 1 && A2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 1) (B2 *> O) = (7.28:7.28:7.28, 9.03:9.03:9.03);
      if (A1 == 0 && A2 == 0 && C1 == 1 && C2 == 0 && D1 == 1 && D2 == 0) (B2 *> O) = (6.73:6.73:6.73, 6.43:6.43:6.43);
      if (A1 == 0 && A2 == 1 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 0) (B2 *> O) = (6.77:6.77:6.77, 7.75:7.75:7.75);
      if (A1 == 0 && A2 == 1 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 1) (B2 *> O) = (6.74:6.74:6.74, 7.75:7.75:7.75);
      if (A1 == 0 && A2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 0) (B2 *> O) = (6.76:6.76:6.76, 6.43:6.43:6.43);
      if (A1 == 0 && A2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 1) (B2 *> O) = (6.73:6.73:6.73, 6.43:6.43:6.43);
      if (A1 == 1 && A2 == 0 && C1 == 0 && C2 == 1 && D1 == 1 && D2 == 0) (B2 *> O) = (7.28:7.28:7.28, 9.03:9.03:9.03);
      if (A1 == 1 && A2 == 0 && C1 == 0 && C2 == 0 && D1 == 1 && D2 == 0) (B2 *> O) = (7.30:7.30:7.30, 9.02:9.02:9.02);
      if (A1 == 1 && A2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 0) (B2 *> O) = (7.31:7.31:7.31, 9.02:9.02:9.02);
      if (A1 == 1 && A2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 0) (B2 *> O) = (7.32:7.32:7.32, 9.01:9.01:9.01);
      if (A1 == 0 && A2 == 1 && C1 == 0 && C2 == 1 && D1 == 1 && D2 == 0) (B2 *> O) = (6.74:6.74:6.74, 7.75:7.75:7.75);
      if (A1 == 1 && A2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 1) (B2 *> O) = (7.28:7.28:7.28, 9.03:9.03:9.03);
      if (A1 == 0 && A2 == 1 && C1 == 0 && C2 == 0 && D1 == 1 && D2 == 0) (B2 *> O) = (6.75:6.75:6.75, 7.75:7.75:7.75);
      if (A1 == 1 && A2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 1) (B2 *> O) = (7.30:7.30:7.30, 9.02:9.02:9.02);
      if (A1 == 0 && A2 == 0 && C1 == 0 && C2 == 1 && D1 == 1 && D2 == 0) (B2 *> O) = (6.73:6.73:6.73, 6.43:6.43:6.43);
      if (A1 == 0 && A2 == 0 && C1 == 0 && C2 == 0 && D1 == 1 && D2 == 0) (B2 *> O) = (6.74:6.74:6.74, 6.43:6.43:6.43);
      if (A1 == 0 && A2 == 1 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 0) (B2 *> O) = (6.77:6.77:6.77, 7.75:7.75:7.75);
      if (A1 == 0 && A2 == 1 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 0) (B2 *> O) = (6.78:6.78:6.78, 7.74:7.74:7.74);
      if (A1 == 0 && A2 == 1 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 1) (B2 *> O) = (6.74:6.74:6.74, 7.75:7.75:7.75);
      if (A1 == 0 && A2 == 1 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 1) (B2 *> O) = (6.75:6.75:6.75, 7.75:7.75:7.75);
      if (A1 == 1 && A2 == 0 && C1 == 1 && C2 == 0 && D1 == 1 && D2 == 0) (B2 *> O) = (7.28:7.28:7.28, 9.03:9.03:9.03);
      if (A1 == 0 && A2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 0) (B2 *> O) = (6.76:6.76:6.76, 6.43:6.43:6.43);
      if (A1 == 0 && A2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 0) (B2 *> O) = (6.77:6.77:6.77, 6.42:6.42:6.42);
      if (A1 == 0 && A2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 1) (B2 *> O) = (6.73:6.73:6.73, 6.43:6.43:6.43);
      ifnone (B2 *> O) = (6.73:6.73:6.73, 6.43:6.43:6.43);
      if (B1 == 1 && B2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 0) (A1 *> O) = (8.19:8.19:8.19, 9.54:9.54:9.54);
      if (B1 == 1 && B2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 0) (A1 *> O) = (8.21:8.21:8.21, 9.53:9.53:9.53);
      if (B1 == 0 && B2 == 1 && C1 == 0 && C2 == 1 && D1 == 1 && D2 == 0) (A1 *> O) = (7.81:7.81:7.81, 8.73:8.73:8.73);
      if (B1 == 1 && B2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 1) (A1 *> O) = (8.17:8.17:8.17, 9.55:9.55:9.55);
      if (B1 == 0 && B2 == 1 && C1 == 0 && C2 == 0 && D1 == 1 && D2 == 0) (A1 *> O) = (7.82:7.82:7.82, 8.73:8.73:8.73);
      if (B1 == 1 && B2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 1) (A1 *> O) = (8.18:8.18:8.18, 9.54:9.54:9.54);
      if (B1 == 0 && B2 == 0 && C1 == 0 && C2 == 1 && D1 == 1 && D2 == 0) (A1 *> O) = (8.15:8.15:8.15, 7.47:7.47:7.47);
      if (B1 == 0 && B2 == 0 && C1 == 0 && C2 == 0 && D1 == 1 && D2 == 0) (A1 *> O) = (8.16:8.16:8.16, 7.47:7.47:7.47);
      if (B1 == 0 && B2 == 1 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 0) (A1 *> O) = (7.83:7.83:7.83, 8.72:8.72:8.72);
      if (B1 == 0 && B2 == 1 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 0) (A1 *> O) = (7.85:7.85:7.85, 8.72:8.72:8.72);
      if (B1 == 0 && B2 == 1 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 1) (A1 *> O) = (7.81:7.81:7.81, 8.73:8.73:8.73);
      if (B1 == 0 && B2 == 1 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 1) (A1 *> O) = (7.82:7.82:7.82, 8.73:8.73:8.73);
      if (B1 == 1 && B2 == 0 && C1 == 1 && C2 == 0 && D1 == 1 && D2 == 0) (A1 *> O) = (8.17:8.17:8.17, 9.55:9.55:9.55);
      if (B1 == 0 && B2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 0) (A1 *> O) = (8.17:8.17:8.17, 7.46:7.46:7.46);
      if (B1 == 0 && B2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 0) (A1 *> O) = (8.19:8.19:8.19, 7.46:7.46:7.46);
      if (B1 == 0 && B2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 1) (A1 *> O) = (8.15:8.15:8.15, 7.47:7.47:7.47);
      if (B1 == 0 && B2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 1) (A1 *> O) = (8.16:8.16:8.16, 7.47:7.47:7.47);
      if (B1 == 1 && B2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 0) (A1 *> O) = (8.19:8.19:8.19, 9.54:9.54:9.54);
      if (B1 == 0 && B2 == 1 && C1 == 1 && C2 == 0 && D1 == 1 && D2 == 0) (A1 *> O) = (7.81:7.81:7.81, 8.73:8.73:8.73);
      if (B1 == 1 && B2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 1) (A1 *> O) = (8.17:8.17:8.17, 9.55:9.55:9.55);
      if (B1 == 0 && B2 == 0 && C1 == 1 && C2 == 0 && D1 == 1 && D2 == 0) (A1 *> O) = (8.15:8.15:8.15, 7.47:7.47:7.47);
      if (B1 == 0 && B2 == 1 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 0) (A1 *> O) = (7.83:7.83:7.83, 8.72:8.72:8.72);
      if (B1 == 0 && B2 == 1 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 1) (A1 *> O) = (7.81:7.81:7.81, 8.73:8.73:8.73);
      if (B1 == 0 && B2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 0) (A1 *> O) = (8.17:8.17:8.17, 7.46:7.46:7.46);
      if (B1 == 0 && B2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 1) (A1 *> O) = (8.15:8.15:8.15, 7.47:7.47:7.47);
      if (B1 == 1 && B2 == 0 && C1 == 0 && C2 == 1 && D1 == 1 && D2 == 0) (A1 *> O) = (8.17:8.17:8.17, 9.55:9.55:9.55);
      if (B1 == 1 && B2 == 0 && C1 == 0 && C2 == 0 && D1 == 1 && D2 == 0) (A1 *> O) = (8.18:8.18:8.18, 9.54:9.54:9.54);
      ifnone (A1 *> O) = (8.18:8.18:8.18, 9.54:9.54:9.54);
      if (B1 == 0 && B2 == 1 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 1) (A2 *> O) = (8.19:8.19:8.19, 9.86:9.86:9.86);
      if (B1 == 0 && B2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 0) (A2 *> O) = (8.55:8.55:8.55, 8.34:8.34:8.34);
      if (B1 == 0 && B2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 1) (A2 *> O) = (8.53:8.53:8.53, 8.35:8.35:8.35);
      if (B1 == 1 && B2 == 0 && C1 == 0 && C2 == 1 && D1 == 1 && D2 == 0) (A2 *> O) = (8.55:8.55:8.55, 10.64:10.64:10.64);
      if (B1 == 1 && B2 == 0 && C1 == 0 && C2 == 0 && D1 == 1 && D2 == 0) (A2 *> O) = (8.56:8.56:8.56, 10.64:10.64:10.64);
      if (B1 == 1 && B2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 0) (A2 *> O) = (8.57:8.57:8.57, 10.64:10.64:10.64);
      if (B1 == 1 && B2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 0) (A2 *> O) = (8.59:8.59:8.59, 10.63:10.63:10.63);
      if (B1 == 1 && B2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 1) (A2 *> O) = (8.55:8.55:8.55, 10.64:10.64:10.64);
      if (B1 == 0 && B2 == 1 && C1 == 0 && C2 == 1 && D1 == 1 && D2 == 0) (A2 *> O) = (8.19:8.19:8.19, 9.86:9.86:9.86);
      if (B1 == 1 && B2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 1) (A2 *> O) = (8.56:8.56:8.56, 10.64:10.64:10.64);
      if (B1 == 0 && B2 == 1 && C1 == 0 && C2 == 0 && D1 == 1 && D2 == 0) (A2 *> O) = (8.20:8.20:8.20, 9.86:9.86:9.86);
      if (B1 == 0 && B2 == 0 && C1 == 0 && C2 == 1 && D1 == 1 && D2 == 0) (A2 *> O) = (8.53:8.53:8.53, 8.35:8.35:8.35);
      if (B1 == 0 && B2 == 0 && C1 == 0 && C2 == 0 && D1 == 1 && D2 == 0) (A2 *> O) = (8.54:8.54:8.54, 8.34:8.34:8.34);
      if (B1 == 0 && B2 == 1 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 0) (A2 *> O) = (8.21:8.21:8.21, 9.85:9.85:9.85);
      if (B1 == 0 && B2 == 1 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 0) (A2 *> O) = (8.23:8.23:8.23, 9.85:9.85:9.85);
      if (B1 == 0 && B2 == 1 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 1) (A2 *> O) = (8.19:8.19:8.19, 9.86:9.86:9.86);
      if (B1 == 0 && B2 == 1 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 1) (A2 *> O) = (8.20:8.20:8.20, 9.86:9.86:9.86);
      if (B1 == 1 && B2 == 0 && C1 == 1 && C2 == 0 && D1 == 1 && D2 == 0) (A2 *> O) = (8.55:8.55:8.55, 10.64:10.64:10.64);
      if (B1 == 0 && B2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 0) (A2 *> O) = (8.55:8.55:8.55, 8.34:8.34:8.34);
      if (B1 == 0 && B2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 0) (A2 *> O) = (8.56:8.56:8.56, 8.34:8.34:8.34);
      if (B1 == 0 && B2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 1) (A2 *> O) = (8.53:8.53:8.53, 8.35:8.35:8.35);
      if (B1 == 0 && B2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 1) (A2 *> O) = (8.54:8.54:8.54, 8.34:8.34:8.34);
      if (B1 == 1 && B2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 0) (A2 *> O) = (8.57:8.57:8.57, 10.64:10.64:10.64);
      if (B1 == 1 && B2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 1) (A2 *> O) = (8.55:8.55:8.55, 10.64:10.64:10.64);
      if (B1 == 0 && B2 == 1 && C1 == 1 && C2 == 0 && D1 == 1 && D2 == 0) (A2 *> O) = (8.19:8.19:8.19, 9.86:9.86:9.86);
      if (B1 == 0 && B2 == 0 && C1 == 1 && C2 == 0 && D1 == 1 && D2 == 0) (A2 *> O) = (8.53:8.53:8.53, 8.35:8.35:8.35);
      if (B1 == 0 && B2 == 1 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 0) (A2 *> O) = (8.21:8.21:8.21, 9.85:9.85:9.85);
      ifnone (A2 *> O) = (8.21:8.21:8.21, 9.85:9.85:9.85);

      //  Module Path Delay
   endspecify
`endprotect
endmodule

`endcelldefine
