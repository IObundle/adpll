// Created by ihdl
`timescale 10ps/1ps

`celldefine

module MAOI1CHD(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;

//Function Block
`protect
   nor g1(o1, B1, B2);
   and g3(o2, A1, A2);
   nor g2(O, o1, o2);

//Specify Block
   specify

      //  Module Path Delay (state dependent)
      if (A1 == 0 && A2 == 1) (B2 *> O) = (5.22:5.22:5.22, 6.23:6.23:6.23);
      if (A1 == 0 && A2 == 0) (B2 *> O) = (4.69:4.69:4.69, 6.22:6.22:6.22);
      if (A1 == 1 && A2 == 0) (B2 *> O) = (6.17:6.17:6.17, 6.37:6.37:6.37);
      ifnone (B2 *> O) = (6.17:6.17:6.17, 6.37:6.37:6.37);
      if (A1 == 1 && A2 == 0) (B1 *> O) = (6.59:6.59:6.59, 7.07:7.07:7.07);
      if (A1 == 0 && A2 == 1) (B1 *> O) = (5.63:5.63:5.63, 6.93:6.93:6.93);
      if (A1 == 0 && A2 == 0) (B1 *> O) = (5.11:5.11:5.11, 6.91:6.91:6.91);
      ifnone (B1 *> O) = (5.11:5.11:5.11, 6.91:6.91:6.91);
      if (B1 == 0 && B2 == 1) (A1 *> O) = (4.78:4.78:4.78, 1.96:1.96:1.96);
      if (B1 == 1 && B2 == 1) (A1 *> O) = (4.73:4.73:4.73, 1.96:1.96:1.96);
      if (B1 == 1 && B2 == 0) (A1 *> O) = (4.78:4.78:4.78, 1.96:1.96:1.96);
      ifnone (A1 *> O) = (4.78:4.78:4.78, 1.96:1.96:1.96);
      if (B1 == 1 && B2 == 0) (A2 *> O) = (5.65:5.65:5.65, 2.04:2.04:2.04);
      if (B1 == 0 && B2 == 1) (A2 *> O) = (5.65:5.65:5.65, 2.04:2.04:2.04);
      if (B1 == 1 && B2 == 1) (A2 *> O) = (5.61:5.61:5.61, 2.04:2.04:2.04);
      ifnone (A2 *> O) = (5.61:5.61:5.61, 2.04:2.04:2.04);

      //  Module Path Delay
   endspecify
`endprotect
endmodule

`endcelldefine
