// Created by ihdl
`timescale 10ps/1ps

`celldefine

module AOI2222KHD(O, A1, A2, B1, B2, C1, C2, D1, D2);
   output O;
   input A1, A2, B1, B2, C1, C2, D1, D2;

//Function Block
`protect
   and g1(o1, B1, B2);
   and g3(o2, A1, A2);
   and g4(o3, C1, C2);
   and g5(o4, D1, D2);
   nor g2(O, o1, o2, o3, o4);

//Specify Block
   specify

      //  Module Path Delay (state dependent)
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 0 && C1 == 0 && C2 == 1) (D1 *> O) = (10.35:10.35:10.35, 8.47:8.47:8.47);
      if (A1 == 1 && A2 == 0 && B1 == 1 && B2 == 0 && C1 == 1 && C2 == 0) (D1 *> O) = (11.93:11.93:11.93, 9.05:9.05:9.05);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 1 && C1 == 0 && C2 == 0) (D1 *> O) = (8.91:8.91:8.91, 8.46:8.46:8.46);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 0 && C1 == 0 && C2 == 0) (D1 *> O) = (8.90:8.90:8.90, 8.46:8.46:8.46);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 1 && C1 == 0 && C2 == 1) (D1 *> O) = (10.35:10.35:10.35, 8.47:8.47:8.47);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 0 && C1 == 0 && C2 == 1) (D1 *> O) = (10.35:10.35:10.35, 8.47:8.47:8.47);
      if (A1 == 1 && A2 == 0 && B1 == 1 && B2 == 0 && C1 == 0 && C2 == 0) (D1 *> O) = (8.91:8.91:8.91, 8.46:8.46:8.46);
      if (A1 == 1 && A2 == 0 && B1 == 1 && B2 == 0 && C1 == 0 && C2 == 1) (D1 *> O) = (10.35:10.35:10.35, 8.47:8.47:8.47);
      if (A1 == 0 && A2 == 1 && B1 == 1 && B2 == 0 && C1 == 1 && C2 == 0) (D1 *> O) = (11.93:11.93:11.93, 9.05:9.05:9.05);
      if (A1 == 0 && A2 == 0 && B1 == 1 && B2 == 0 && C1 == 1 && C2 == 0) (D1 *> O) = (11.93:11.93:11.93, 9.06:9.06:9.06);
      if (A1 == 0 && A2 == 1 && B1 == 1 && B2 == 0 && C1 == 0 && C2 == 0) (D1 *> O) = (8.91:8.91:8.91, 8.46:8.46:8.46);
      if (A1 == 0 && A2 == 1 && B1 == 1 && B2 == 0 && C1 == 0 && C2 == 1) (D1 *> O) = (10.35:10.35:10.35, 8.47:8.47:8.47);
      if (A1 == 0 && A2 == 0 && B1 == 1 && B2 == 0 && C1 == 0 && C2 == 0) (D1 *> O) = (8.91:8.91:8.91, 8.46:8.46:8.46);
      if (A1 == 0 && A2 == 0 && B1 == 1 && B2 == 0 && C1 == 0 && C2 == 1) (D1 *> O) = (10.35:10.35:10.35, 8.47:8.47:8.47);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 1 && C1 == 1 && C2 == 0) (D1 *> O) = (11.93:11.93:11.93, 9.05:9.05:9.05);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 0 && C1 == 1 && C2 == 0) (D1 *> O) = (11.93:11.93:11.93, 9.06:9.06:9.06);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 1 && C1 == 0 && C2 == 0) (D1 *> O) = (8.91:8.91:8.91, 8.46:8.46:8.46);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 0 && C1 == 0 && C2 == 0) (D1 *> O) = (8.90:8.90:8.90, 8.46:8.46:8.46);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 1 && C1 == 0 && C2 == 1) (D1 *> O) = (10.35:10.35:10.35, 8.47:8.47:8.47);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 1 && C1 == 1 && C2 == 0) (D1 *> O) = (11.93:11.93:11.93, 9.05:9.05:9.05);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 0 && C1 == 0 && C2 == 1) (D1 *> O) = (10.35:10.35:10.35, 8.47:8.47:8.47);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 0 && C1 == 1 && C2 == 0) (D1 *> O) = (11.93:11.93:11.93, 9.06:9.06:9.06);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 1 && C1 == 1 && C2 == 0) (D1 *> O) = (11.93:11.93:11.93, 9.06:9.06:9.06);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 0 && C1 == 1 && C2 == 0) (D1 *> O) = (11.93:11.93:11.93, 9.06:9.06:9.06);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 1 && C1 == 0 && C2 == 0) (D1 *> O) = (8.91:8.91:8.91, 8.46:8.46:8.46);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 0 && C1 == 0 && C2 == 0) (D1 *> O) = (8.90:8.90:8.90, 8.46:8.46:8.46);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 1 && C1 == 0 && C2 == 1) (D1 *> O) = (10.35:10.35:10.35, 8.47:8.47:8.47);
      ifnone (D1 *> O) = (10.35:10.35:10.35, 8.47:8.47:8.47);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 1 && C1 == 1 && C2 == 0) (D2 *> O) = (12.70:12.70:12.70, 9.13:9.13:9.13);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 0 && C1 == 1 && C2 == 0) (D2 *> O) = (12.70:12.70:12.70, 9.13:9.13:9.13);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 1 && C1 == 0 && C2 == 0) (D2 *> O) = (9.50:9.50:9.50, 8.53:8.53:8.53);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 0 && C1 == 0 && C2 == 0) (D2 *> O) = (9.50:9.50:9.50, 8.53:8.53:8.53);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 1 && C1 == 1 && C2 == 0) (D2 *> O) = (12.70:12.70:12.70, 9.13:9.13:9.13);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 1 && C1 == 0 && C2 == 1) (D2 *> O) = (11.14:11.14:11.14, 8.54:8.54:8.54);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 0 && C1 == 0 && C2 == 1) (D2 *> O) = (11.14:11.14:11.14, 8.54:8.54:8.54);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 0 && C1 == 1 && C2 == 0) (D2 *> O) = (12.70:12.70:12.70, 9.13:9.13:9.13);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 1 && C1 == 1 && C2 == 0) (D2 *> O) = (12.70:12.70:12.70, 9.13:9.13:9.13);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 0 && C1 == 1 && C2 == 0) (D2 *> O) = (12.70:12.70:12.70, 9.13:9.13:9.13);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 1 && C1 == 0 && C2 == 0) (D2 *> O) = (9.50:9.50:9.50, 8.53:8.53:8.53);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 0 && C1 == 0 && C2 == 0) (D2 *> O) = (9.50:9.50:9.50, 8.53:8.53:8.53);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 1 && C1 == 0 && C2 == 1) (D2 *> O) = (11.14:11.14:11.14, 8.54:8.54:8.54);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 0 && C1 == 0 && C2 == 1) (D2 *> O) = (11.14:11.14:11.14, 8.54:8.54:8.54);
      if (A1 == 1 && A2 == 0 && B1 == 1 && B2 == 0 && C1 == 1 && C2 == 0) (D2 *> O) = (12.70:12.70:12.70, 9.13:9.13:9.13);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 1 && C1 == 0 && C2 == 0) (D2 *> O) = (9.50:9.50:9.50, 8.53:8.53:8.53);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 0 && C1 == 0 && C2 == 0) (D2 *> O) = (9.50:9.50:9.50, 8.54:8.54:8.54);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 1 && C1 == 0 && C2 == 1) (D2 *> O) = (11.14:11.14:11.14, 8.54:8.54:8.54);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 0 && C1 == 0 && C2 == 1) (D2 *> O) = (11.14:11.14:11.14, 8.54:8.54:8.54);
      if (A1 == 1 && A2 == 0 && B1 == 1 && B2 == 0 && C1 == 0 && C2 == 0) (D2 *> O) = (9.50:9.50:9.50, 8.53:8.53:8.53);
      if (A1 == 0 && A2 == 1 && B1 == 1 && B2 == 0 && C1 == 1 && C2 == 0) (D2 *> O) = (12.70:12.70:12.70, 9.13:9.13:9.13);
      if (A1 == 1 && A2 == 0 && B1 == 1 && B2 == 0 && C1 == 0 && C2 == 1) (D2 *> O) = (11.14:11.14:11.14, 8.54:8.54:8.54);
      if (A1 == 0 && A2 == 0 && B1 == 1 && B2 == 0 && C1 == 1 && C2 == 0) (D2 *> O) = (12.70:12.70:12.70, 9.13:9.13:9.13);
      if (A1 == 0 && A2 == 1 && B1 == 1 && B2 == 0 && C1 == 0 && C2 == 0) (D2 *> O) = (9.50:9.50:9.50, 8.53:8.53:8.53);
      if (A1 == 0 && A2 == 1 && B1 == 1 && B2 == 0 && C1 == 0 && C2 == 1) (D2 *> O) = (11.14:11.14:11.14, 8.54:8.54:8.54);
      if (A1 == 0 && A2 == 0 && B1 == 1 && B2 == 0 && C1 == 0 && C2 == 0) (D2 *> O) = (9.50:9.50:9.50, 8.53:8.53:8.53);
      if (A1 == 0 && A2 == 0 && B1 == 1 && B2 == 0 && C1 == 0 && C2 == 1) (D2 *> O) = (11.14:11.14:11.14, 8.54:8.54:8.54);
      ifnone (D2 *> O) = (11.14:11.14:11.14, 8.54:8.54:8.54);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 0 && D1 == 0 && D2 == 0) (C1 *> O) = (10.62:10.62:10.62, 9.65:9.65:9.65);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 1 && D1 == 0 && D2 == 1) (C1 *> O) = (12.03:12.03:12.03, 9.34:9.34:9.34);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 0 && D1 == 0 && D2 == 1) (C1 *> O) = (12.03:12.03:12.03, 9.34:9.34:9.34);
      if (A1 == 1 && A2 == 0 && B1 == 1 && B2 == 0 && D1 == 1 && D2 == 0) (C1 *> O) = (12.96:12.96:12.96, 9.68:9.68:9.68);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 1 && D1 == 0 && D2 == 0) (C1 *> O) = (10.62:10.62:10.62, 9.65:9.65:9.65);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 0 && D1 == 0 && D2 == 0) (C1 *> O) = (10.62:10.62:10.62, 9.65:9.65:9.65);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 1 && D1 == 0 && D2 == 1) (C1 *> O) = (12.03:12.03:12.03, 9.34:9.34:9.34);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 0 && D1 == 0 && D2 == 1) (C1 *> O) = (12.03:12.03:12.03, 9.34:9.34:9.34);
      if (A1 == 1 && A2 == 0 && B1 == 1 && B2 == 0 && D1 == 0 && D2 == 0) (C1 *> O) = (10.62:10.62:10.62, 9.65:9.65:9.65);
      if (A1 == 0 && A2 == 1 && B1 == 1 && B2 == 0 && D1 == 1 && D2 == 0) (C1 *> O) = (12.96:12.96:12.96, 9.68:9.68:9.68);
      if (A1 == 1 && A2 == 0 && B1 == 1 && B2 == 0 && D1 == 0 && D2 == 1) (C1 *> O) = (12.03:12.03:12.03, 9.34:9.34:9.34);
      if (A1 == 0 && A2 == 0 && B1 == 1 && B2 == 0 && D1 == 1 && D2 == 0) (C1 *> O) = (12.96:12.96:12.96, 9.68:9.68:9.68);
      if (A1 == 0 && A2 == 1 && B1 == 1 && B2 == 0 && D1 == 0 && D2 == 0) (C1 *> O) = (10.62:10.62:10.62, 9.65:9.65:9.65);
      if (A1 == 0 && A2 == 1 && B1 == 1 && B2 == 0 && D1 == 0 && D2 == 1) (C1 *> O) = (12.03:12.03:12.03, 9.34:9.34:9.34);
      if (A1 == 0 && A2 == 0 && B1 == 1 && B2 == 0 && D1 == 0 && D2 == 0) (C1 *> O) = (10.62:10.62:10.62, 9.65:9.65:9.65);
      if (A1 == 0 && A2 == 0 && B1 == 1 && B2 == 0 && D1 == 0 && D2 == 1) (C1 *> O) = (12.03:12.03:12.03, 9.34:9.34:9.34);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 1 && D1 == 1 && D2 == 0) (C1 *> O) = (12.96:12.96:12.96, 9.68:9.68:9.68);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 0 && D1 == 1 && D2 == 0) (C1 *> O) = (12.96:12.96:12.96, 9.68:9.68:9.68);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 1 && D1 == 0 && D2 == 0) (C1 *> O) = (10.62:10.62:10.62, 9.65:9.65:9.65);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 0 && D1 == 0 && D2 == 0) (C1 *> O) = (10.62:10.62:10.62, 9.65:9.65:9.65);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 1 && D1 == 1 && D2 == 0) (C1 *> O) = (12.96:12.96:12.96, 9.68:9.68:9.68);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 1 && D1 == 0 && D2 == 1) (C1 *> O) = (12.03:12.03:12.03, 9.34:9.34:9.34);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 0 && D1 == 1 && D2 == 0) (C1 *> O) = (12.96:12.96:12.96, 9.68:9.68:9.68);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 0 && D1 == 0 && D2 == 1) (C1 *> O) = (12.03:12.03:12.03, 9.34:9.34:9.34);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 1 && D1 == 1 && D2 == 0) (C1 *> O) = (12.96:12.96:12.96, 9.68:9.68:9.68);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 0 && D1 == 1 && D2 == 0) (C1 *> O) = (12.96:12.96:12.96, 9.68:9.68:9.68);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 1 && D1 == 0 && D2 == 0) (C1 *> O) = (10.62:10.62:10.62, 9.65:9.65:9.65);
      ifnone (C1 *> O) = (10.62:10.62:10.62, 9.65:9.65:9.65);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 1 && D1 == 1 && D2 == 0) (C2 *> O) = (14.39:14.39:14.39, 10.00:10.00:10.00);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 0 && D1 == 1 && D2 == 0) (C2 *> O) = (14.39:14.39:14.39, 10.00:10.00:10.00);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 1 && D1 == 0 && D2 == 0) (C2 *> O) = (11.72:11.72:11.72, 9.97:9.97:9.97);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 0 && D1 == 0 && D2 == 0) (C2 *> O) = (11.72:11.72:11.72, 9.97:9.97:9.97);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 1 && D1 == 1 && D2 == 0) (C2 *> O) = (14.39:14.39:14.39, 10.00:10.00:10.00);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 1 && D1 == 0 && D2 == 1) (C2 *> O) = (13.47:13.47:13.47, 9.66:9.66:9.66);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 0 && D1 == 1 && D2 == 0) (C2 *> O) = (14.39:14.39:14.39, 10.00:10.00:10.00);
      if (A1 == 1 && A2 == 0 && B1 == 0 && B2 == 0 && D1 == 0 && D2 == 1) (C2 *> O) = (13.47:13.47:13.47, 9.66:9.66:9.66);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 1 && D1 == 1 && D2 == 0) (C2 *> O) = (14.39:14.39:14.39, 10.00:10.00:10.00);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 0 && D1 == 1 && D2 == 0) (C2 *> O) = (14.39:14.39:14.39, 10.00:10.00:10.00);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 1 && D1 == 0 && D2 == 0) (C2 *> O) = (11.72:11.72:11.72, 9.97:9.97:9.97);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 0 && D1 == 0 && D2 == 0) (C2 *> O) = (11.72:11.72:11.72, 9.97:9.97:9.97);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 1 && D1 == 0 && D2 == 1) (C2 *> O) = (13.47:13.47:13.47, 9.66:9.66:9.66);
      if (A1 == 0 && A2 == 1 && B1 == 0 && B2 == 0 && D1 == 0 && D2 == 1) (C2 *> O) = (13.47:13.47:13.47, 9.66:9.66:9.66);
      if (A1 == 1 && A2 == 0 && B1 == 1 && B2 == 0 && D1 == 1 && D2 == 0) (C2 *> O) = (14.39:14.39:14.39, 10.00:10.00:10.00);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 1 && D1 == 0 && D2 == 0) (C2 *> O) = (11.72:11.72:11.72, 9.97:9.97:9.97);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 0 && D1 == 0 && D2 == 0) (C2 *> O) = (11.72:11.72:11.72, 9.97:9.97:9.97);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 1 && D1 == 0 && D2 == 1) (C2 *> O) = (13.47:13.47:13.47, 9.66:9.66:9.66);
      if (A1 == 0 && A2 == 0 && B1 == 0 && B2 == 0 && D1 == 0 && D2 == 1) (C2 *> O) = (13.47:13.47:13.47, 9.66:9.66:9.66);
      if (A1 == 1 && A2 == 0 && B1 == 1 && B2 == 0 && D1 == 0 && D2 == 0) (C2 *> O) = (11.72:11.72:11.72, 9.97:9.97:9.97);
      if (A1 == 0 && A2 == 1 && B1 == 1 && B2 == 0 && D1 == 1 && D2 == 0) (C2 *> O) = (14.39:14.39:14.39, 10.00:10.00:10.00);
      if (A1 == 1 && A2 == 0 && B1 == 1 && B2 == 0 && D1 == 0 && D2 == 1) (C2 *> O) = (13.47:13.47:13.47, 9.66:9.66:9.66);
      if (A1 == 0 && A2 == 0 && B1 == 1 && B2 == 0 && D1 == 1 && D2 == 0) (C2 *> O) = (14.39:14.39:14.39, 10.00:10.00:10.00);
      if (A1 == 0 && A2 == 1 && B1 == 1 && B2 == 0 && D1 == 0 && D2 == 0) (C2 *> O) = (11.72:11.72:11.72, 9.97:9.97:9.97);
      if (A1 == 0 && A2 == 1 && B1 == 1 && B2 == 0 && D1 == 0 && D2 == 1) (C2 *> O) = (13.47:13.47:13.47, 9.66:9.66:9.66);
      if (A1 == 0 && A2 == 0 && B1 == 1 && B2 == 0 && D1 == 0 && D2 == 0) (C2 *> O) = (11.72:11.72:11.72, 9.97:9.97:9.97);
      if (A1 == 0 && A2 == 0 && B1 == 1 && B2 == 0 && D1 == 0 && D2 == 1) (C2 *> O) = (13.47:13.47:13.47, 9.66:9.66:9.66);
      ifnone (C2 *> O) = (13.47:13.47:13.47, 9.66:9.66:9.66);
      if (A1 == 1 && A2 == 0 && C1 == 0 && C2 == 1 && D1 == 1 && D2 == 0) (B1 *> O) = (11.96:11.96:11.96, 9.67:9.67:9.67);
      if (A1 == 1 && A2 == 0 && C1 == 0 && C2 == 0 && D1 == 1 && D2 == 0) (B1 *> O) = (11.95:11.95:11.95, 9.68:9.68:9.68);
      if (A1 == 1 && A2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 0) (B1 *> O) = (11.95:11.95:11.95, 9.69:9.69:9.69);
      if (A1 == 1 && A2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 0) (B1 *> O) = (11.93:11.93:11.93, 9.70:9.70:9.70);
      if (A1 == 0 && A2 == 1 && C1 == 0 && C2 == 1 && D1 == 1 && D2 == 0) (B1 *> O) = (10.50:10.50:10.50, 9.10:9.10:9.10);
      if (A1 == 1 && A2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 1) (B1 *> O) = (11.96:11.96:11.96, 9.67:9.67:9.67);
      if (A1 == 0 && A2 == 1 && C1 == 0 && C2 == 0 && D1 == 1 && D2 == 0) (B1 *> O) = (10.49:10.49:10.49, 9.11:9.11:9.11);
      if (A1 == 1 && A2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 1) (B1 *> O) = (11.95:11.95:11.95, 9.68:9.68:9.68);
      if (A1 == 0 && A2 == 0 && C1 == 0 && C2 == 1 && D1 == 1 && D2 == 0) (B1 *> O) = (9.08:9.08:9.08, 9.09:9.09:9.09);
      if (A1 == 0 && A2 == 0 && C1 == 0 && C2 == 0 && D1 == 1 && D2 == 0) (B1 *> O) = (9.07:9.07:9.07, 9.10:9.10:9.10);
      if (A1 == 0 && A2 == 1 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 0) (B1 *> O) = (10.48:10.48:10.48, 9.12:9.12:9.12);
      if (A1 == 0 && A2 == 1 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 0) (B1 *> O) = (10.47:10.47:10.47, 9.13:9.13:9.13);
      if (A1 == 0 && A2 == 1 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 1) (B1 *> O) = (10.50:10.50:10.50, 9.10:9.10:9.10);
      if (A1 == 0 && A2 == 1 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 1) (B1 *> O) = (10.49:10.49:10.49, 9.11:9.11:9.11);
      if (A1 == 1 && A2 == 0 && C1 == 1 && C2 == 0 && D1 == 1 && D2 == 0) (B1 *> O) = (11.96:11.96:11.96, 9.67:9.67:9.67);
      if (A1 == 0 && A2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 0) (B1 *> O) = (9.05:9.05:9.05, 9.11:9.11:9.11);
      if (A1 == 0 && A2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 0) (B1 *> O) = (9.04:9.04:9.04, 9.12:9.12:9.12);
      if (A1 == 0 && A2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 1) (B1 *> O) = (9.08:9.08:9.08, 9.09:9.09:9.09);
      if (A1 == 0 && A2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 1) (B1 *> O) = (9.07:9.07:9.07, 9.10:9.10:9.10);
      if (A1 == 1 && A2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 0) (B1 *> O) = (11.95:11.95:11.95, 9.69:9.69:9.69);
      if (A1 == 0 && A2 == 1 && C1 == 1 && C2 == 0 && D1 == 1 && D2 == 0) (B1 *> O) = (10.50:10.50:10.50, 9.10:9.10:9.10);
      if (A1 == 1 && A2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 1) (B1 *> O) = (11.96:11.96:11.96, 9.67:9.67:9.67);
      if (A1 == 0 && A2 == 0 && C1 == 1 && C2 == 0 && D1 == 1 && D2 == 0) (B1 *> O) = (9.08:9.08:9.08, 9.09:9.09:9.09);
      if (A1 == 0 && A2 == 1 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 0) (B1 *> O) = (10.48:10.48:10.48, 9.12:9.12:9.12);
      if (A1 == 0 && A2 == 1 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 1) (B1 *> O) = (10.50:10.50:10.50, 9.10:9.10:9.10);
      if (A1 == 0 && A2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 0) (B1 *> O) = (9.05:9.05:9.05, 9.11:9.11:9.11);
      if (A1 == 0 && A2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 1) (B1 *> O) = (9.08:9.08:9.08, 9.09:9.09:9.09);
      ifnone (B1 *> O) = (9.08:9.08:9.08, 9.09:9.09:9.09);
      if (A1 == 0 && A2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 1) (B2 *> O) = (9.64:9.64:9.64, 9.18:9.18:9.18);
      if (A1 == 1 && A2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 0) (B2 *> O) = (12.70:12.70:12.70, 9.76:9.76:9.76);
      if (A1 == 0 && A2 == 1 && C1 == 1 && C2 == 0 && D1 == 1 && D2 == 0) (B2 *> O) = (11.27:11.27:11.27, 9.18:9.18:9.18);
      if (A1 == 1 && A2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 1) (B2 *> O) = (12.71:12.71:12.71, 9.74:9.74:9.74);
      if (A1 == 0 && A2 == 0 && C1 == 1 && C2 == 0 && D1 == 1 && D2 == 0) (B2 *> O) = (9.65:9.65:9.65, 9.17:9.17:9.17);
      if (A1 == 0 && A2 == 1 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 0) (B2 *> O) = (11.25:11.25:11.25, 9.19:9.19:9.19);
      if (A1 == 0 && A2 == 1 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 1) (B2 *> O) = (11.27:11.27:11.27, 9.18:9.18:9.18);
      if (A1 == 0 && A2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 0) (B2 *> O) = (9.63:9.63:9.63, 9.18:9.18:9.18);
      if (A1 == 0 && A2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 1) (B2 *> O) = (9.65:9.65:9.65, 9.17:9.17:9.17);
      if (A1 == 1 && A2 == 0 && C1 == 0 && C2 == 1 && D1 == 1 && D2 == 0) (B2 *> O) = (12.71:12.71:12.71, 9.74:9.74:9.74);
      if (A1 == 1 && A2 == 0 && C1 == 0 && C2 == 0 && D1 == 1 && D2 == 0) (B2 *> O) = (12.70:12.70:12.70, 9.75:9.75:9.75);
      if (A1 == 1 && A2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 0) (B2 *> O) = (12.70:12.70:12.70, 9.76:9.76:9.76);
      if (A1 == 1 && A2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 0) (B2 *> O) = (12.69:12.69:12.69, 9.77:9.77:9.77);
      if (A1 == 0 && A2 == 1 && C1 == 0 && C2 == 1 && D1 == 1 && D2 == 0) (B2 *> O) = (11.27:11.27:11.27, 9.18:9.18:9.18);
      if (A1 == 1 && A2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 1) (B2 *> O) = (12.71:12.71:12.71, 9.74:9.74:9.74);
      if (A1 == 0 && A2 == 1 && C1 == 0 && C2 == 0 && D1 == 1 && D2 == 0) (B2 *> O) = (11.26:11.26:11.26, 9.19:9.19:9.19);
      if (A1 == 1 && A2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 1) (B2 *> O) = (12.70:12.70:12.70, 9.75:9.75:9.75);
      if (A1 == 0 && A2 == 0 && C1 == 0 && C2 == 1 && D1 == 1 && D2 == 0) (B2 *> O) = (9.65:9.65:9.65, 9.17:9.17:9.17);
      if (A1 == 0 && A2 == 0 && C1 == 0 && C2 == 0 && D1 == 1 && D2 == 0) (B2 *> O) = (9.64:9.64:9.64, 9.18:9.18:9.18);
      if (A1 == 0 && A2 == 1 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 0) (B2 *> O) = (11.25:11.25:11.25, 9.19:9.19:9.19);
      if (A1 == 0 && A2 == 1 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 0) (B2 *> O) = (11.24:11.24:11.24, 9.20:9.20:9.20);
      if (A1 == 0 && A2 == 1 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 1) (B2 *> O) = (11.27:11.27:11.27, 9.18:9.18:9.18);
      if (A1 == 0 && A2 == 1 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 1) (B2 *> O) = (11.26:11.26:11.26, 9.19:9.19:9.19);
      if (A1 == 1 && A2 == 0 && C1 == 1 && C2 == 0 && D1 == 1 && D2 == 0) (B2 *> O) = (12.71:12.71:12.71, 9.74:9.74:9.74);
      if (A1 == 0 && A2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 0) (B2 *> O) = (9.63:9.63:9.63, 9.18:9.18:9.18);
      if (A1 == 0 && A2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 0) (B2 *> O) = (9.62:9.62:9.62, 9.19:9.19:9.19);
      if (A1 == 0 && A2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 1) (B2 *> O) = (9.65:9.65:9.65, 9.17:9.17:9.17);
      ifnone (B2 *> O) = (9.65:9.65:9.65, 9.17:9.17:9.17);
      if (B1 == 1 && B2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 0) (A1 *> O) = (13.04:13.04:13.04, 10.66:10.66:10.66);
      if (B1 == 1 && B2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 0) (A1 *> O) = (13.03:13.03:13.03, 10.67:10.67:10.67);
      if (B1 == 0 && B2 == 1 && C1 == 0 && C2 == 1 && D1 == 1 && D2 == 0) (A1 *> O) = (12.15:12.15:12.15, 10.28:10.28:10.28);
      if (B1 == 1 && B2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 1) (A1 *> O) = (13.06:13.06:13.06, 10.65:10.65:10.65);
      if (B1 == 0 && B2 == 1 && C1 == 0 && C2 == 0 && D1 == 1 && D2 == 0) (A1 *> O) = (12.14:12.14:12.14, 10.29:10.29:10.29);
      if (B1 == 1 && B2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 1) (A1 *> O) = (13.05:13.05:13.05, 10.66:10.66:10.66);
      if (B1 == 0 && B2 == 0 && C1 == 0 && C2 == 1 && D1 == 1 && D2 == 0) (A1 *> O) = (10.73:10.73:10.73, 10.60:10.60:10.60);
      if (B1 == 0 && B2 == 0 && C1 == 0 && C2 == 0 && D1 == 1 && D2 == 0) (A1 *> O) = (10.72:10.72:10.72, 10.61:10.61:10.61);
      if (B1 == 0 && B2 == 1 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 0) (A1 *> O) = (12.13:12.13:12.13, 10.29:10.29:10.29);
      if (B1 == 0 && B2 == 1 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 0) (A1 *> O) = (12.12:12.12:12.12, 10.30:10.30:10.30);
      if (B1 == 0 && B2 == 1 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 1) (A1 *> O) = (12.15:12.15:12.15, 10.28:10.28:10.28);
      if (B1 == 0 && B2 == 1 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 1) (A1 *> O) = (12.14:12.14:12.14, 10.29:10.29:10.29);
      if (B1 == 1 && B2 == 0 && C1 == 1 && C2 == 0 && D1 == 1 && D2 == 0) (A1 *> O) = (13.06:13.06:13.06, 10.65:10.65:10.65);
      if (B1 == 0 && B2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 0) (A1 *> O) = (10.70:10.70:10.70, 10.62:10.62:10.62);
      if (B1 == 0 && B2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 0) (A1 *> O) = (10.69:10.69:10.69, 10.63:10.63:10.63);
      if (B1 == 0 && B2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 1) (A1 *> O) = (10.73:10.73:10.73, 10.60:10.60:10.60);
      if (B1 == 0 && B2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 1) (A1 *> O) = (10.72:10.72:10.72, 10.61:10.61:10.61);
      if (B1 == 1 && B2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 0) (A1 *> O) = (13.04:13.04:13.04, 10.66:10.66:10.66);
      if (B1 == 0 && B2 == 1 && C1 == 1 && C2 == 0 && D1 == 1 && D2 == 0) (A1 *> O) = (12.15:12.15:12.15, 10.28:10.28:10.28);
      if (B1 == 1 && B2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 1) (A1 *> O) = (13.06:13.06:13.06, 10.65:10.65:10.65);
      if (B1 == 0 && B2 == 0 && C1 == 1 && C2 == 0 && D1 == 1 && D2 == 0) (A1 *> O) = (10.73:10.73:10.73, 10.60:10.60:10.60);
      if (B1 == 0 && B2 == 1 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 0) (A1 *> O) = (12.13:12.13:12.13, 10.29:10.29:10.29);
      if (B1 == 0 && B2 == 1 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 1) (A1 *> O) = (12.15:12.15:12.15, 10.28:10.28:10.28);
      if (B1 == 0 && B2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 0) (A1 *> O) = (10.70:10.70:10.70, 10.62:10.62:10.62);
      if (B1 == 0 && B2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 1) (A1 *> O) = (10.73:10.73:10.73, 10.60:10.60:10.60);
      if (B1 == 1 && B2 == 0 && C1 == 0 && C2 == 1 && D1 == 1 && D2 == 0) (A1 *> O) = (13.06:13.06:13.06, 10.65:10.65:10.65);
      if (B1 == 1 && B2 == 0 && C1 == 0 && C2 == 0 && D1 == 1 && D2 == 0) (A1 *> O) = (13.05:13.05:13.05, 10.66:10.66:10.66);
      ifnone (A1 *> O) = (13.05:13.05:13.05, 10.66:10.66:10.66);
      if (B1 == 0 && B2 == 1 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 1) (A2 *> O) = (13.43:13.43:13.43, 10.65:10.65:10.65);
      if (B1 == 0 && B2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 0) (A2 *> O) = (11.69:11.69:11.69, 10.99:10.99:10.99);
      if (B1 == 0 && B2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 1) (A2 *> O) = (11.71:11.71:11.71, 10.98:10.98:10.98);
      if (B1 == 1 && B2 == 0 && C1 == 0 && C2 == 1 && D1 == 1 && D2 == 0) (A2 *> O) = (14.33:14.33:14.33, 11.03:11.03:11.03);
      if (B1 == 1 && B2 == 0 && C1 == 0 && C2 == 0 && D1 == 1 && D2 == 0) (A2 *> O) = (14.32:14.32:14.32, 11.04:11.04:11.04);
      if (B1 == 1 && B2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 0) (A2 *> O) = (14.31:14.31:14.31, 11.04:11.04:11.04);
      if (B1 == 1 && B2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 0) (A2 *> O) = (14.30:14.30:14.30, 11.05:11.05:11.05);
      if (B1 == 1 && B2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 1) (A2 *> O) = (14.33:14.33:14.33, 11.03:11.03:11.03);
      if (B1 == 0 && B2 == 1 && C1 == 0 && C2 == 1 && D1 == 1 && D2 == 0) (A2 *> O) = (13.43:13.43:13.43, 10.65:10.65:10.65);
      if (B1 == 1 && B2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 1) (A2 *> O) = (14.32:14.32:14.32, 11.04:11.04:11.04);
      if (B1 == 0 && B2 == 1 && C1 == 0 && C2 == 0 && D1 == 1 && D2 == 0) (A2 *> O) = (13.42:13.42:13.42, 10.66:10.66:10.66);
      if (B1 == 0 && B2 == 0 && C1 == 0 && C2 == 1 && D1 == 1 && D2 == 0) (A2 *> O) = (11.71:11.71:11.71, 10.98:10.98:10.98);
      if (B1 == 0 && B2 == 0 && C1 == 0 && C2 == 0 && D1 == 1 && D2 == 0) (A2 *> O) = (11.70:11.70:11.70, 10.99:10.99:10.99);
      if (B1 == 0 && B2 == 1 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 0) (A2 *> O) = (13.41:13.41:13.41, 10.67:10.67:10.67);
      if (B1 == 0 && B2 == 1 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 0) (A2 *> O) = (13.40:13.40:13.40, 10.68:10.68:10.68);
      if (B1 == 0 && B2 == 1 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 1) (A2 *> O) = (13.43:13.43:13.43, 10.65:10.65:10.65);
      if (B1 == 0 && B2 == 1 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 1) (A2 *> O) = (13.42:13.42:13.42, 10.66:10.66:10.66);
      if (B1 == 1 && B2 == 0 && C1 == 1 && C2 == 0 && D1 == 1 && D2 == 0) (A2 *> O) = (14.33:14.33:14.33, 11.03:11.03:11.03);
      if (B1 == 0 && B2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 0) (A2 *> O) = (11.69:11.69:11.69, 10.99:10.99:10.99);
      if (B1 == 0 && B2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 0) (A2 *> O) = (11.68:11.68:11.68, 11.01:11.01:11.01);
      if (B1 == 0 && B2 == 0 && C1 == 0 && C2 == 1 && D1 == 0 && D2 == 1) (A2 *> O) = (11.71:11.71:11.71, 10.98:10.98:10.98);
      if (B1 == 0 && B2 == 0 && C1 == 0 && C2 == 0 && D1 == 0 && D2 == 1) (A2 *> O) = (11.70:11.70:11.70, 10.99:10.99:10.99);
      if (B1 == 1 && B2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 0) (A2 *> O) = (14.31:14.31:14.31, 11.04:11.04:11.04);
      if (B1 == 1 && B2 == 0 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 1) (A2 *> O) = (14.33:14.33:14.33, 11.03:11.03:11.03);
      if (B1 == 0 && B2 == 1 && C1 == 1 && C2 == 0 && D1 == 1 && D2 == 0) (A2 *> O) = (13.43:13.43:13.43, 10.65:10.65:10.65);
      if (B1 == 0 && B2 == 0 && C1 == 1 && C2 == 0 && D1 == 1 && D2 == 0) (A2 *> O) = (11.71:11.71:11.71, 10.98:10.98:10.98);
      if (B1 == 0 && B2 == 1 && C1 == 1 && C2 == 0 && D1 == 0 && D2 == 0) (A2 *> O) = (13.41:13.41:13.41, 10.67:10.67:10.67);
      ifnone (A2 *> O) = (13.41:13.41:13.41, 10.67:10.67:10.67);

      //  Module Path Delay
   endspecify
`endprotect
endmodule

`endcelldefine
