// Created by ihdl
`timescale 10ps/1ps

`celldefine

module MAOI1HHD(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;

//Function Block
`protect
   nor g1(o1, B1, B2);
   and g3(o2, A1, A2);
   nor g2(O, o1, o2);

//Specify Block
   specify

      //  Module Path Delay (state dependent)
      if (A1 == 0 && A2 == 1) (B2 *> O) = (5.07:5.07:5.07, 7.15:7.15:7.15);
      if (A1 == 0 && A2 == 0) (B2 *> O) = (5.07:5.07:5.07, 7.16:7.16:7.16);
      if (A1 == 1 && A2 == 0) (B2 *> O) = (5.07:5.07:5.07, 7.15:7.15:7.15);
      ifnone (B2 *> O) = (5.07:5.07:5.07, 7.15:7.15:7.15);
      if (A1 == 1 && A2 == 0) (B1 *> O) = (4.57:4.57:4.57, 6.49:6.49:6.49);
      if (A1 == 0 && A2 == 1) (B1 *> O) = (4.57:4.57:4.57, 6.49:6.49:6.49);
      if (A1 == 0 && A2 == 0) (B1 *> O) = (4.57:4.57:4.57, 6.49:6.49:6.49);
      ifnone (B1 *> O) = (4.57:4.57:4.57, 6.49:6.49:6.49);
      if (B1 == 0 && B2 == 1) (A1 *> O) = (9.42:9.42:9.42, 8.82:8.82:8.82);
      if (B1 == 1 && B2 == 1) (A1 *> O) = (8.44:8.44:8.44, 8.90:8.90:8.90);
      if (B1 == 1 && B2 == 0) (A1 *> O) = (8.82:8.82:8.82, 8.66:8.66:8.66);
      ifnone (A1 *> O) = (8.82:8.82:8.82, 8.66:8.66:8.66);
      if (B1 == 1 && B2 == 0) (A2 *> O) = (9.36:9.36:9.36, 8.74:8.74:8.74);
      if (B1 == 0 && B2 == 1) (A2 *> O) = (9.97:9.97:9.97, 8.91:8.91:8.91);
      if (B1 == 1 && B2 == 1) (A2 *> O) = (8.99:8.99:8.99, 8.99:8.99:8.99);
      ifnone (A2 *> O) = (8.99:8.99:8.99, 8.99:8.99:8.99);

      //  Module Path Delay
   endspecify
`endprotect
endmodule

`endcelldefine
